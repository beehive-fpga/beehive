`ifndef UDP_RS_ENCODE_DEFS_SVH
`define UDP_RS_ENCODE_DEFS_SVH
    `include "noc_defs.vh"
    `include "packet_defs.vh"

    import udp_rs_encode_pkg::*;

    import beehive_udp_msg::*;
    import beehive_rs_app_stats_msg::*;

`endif
