`ifndef UDP_ECHO_APP_STATS_DEFS_SVH
`define UDP_ECHO_APP_STATS_DEFS_SVH

    `include "noc_defs.vh"

    import beehive_noc_msg::*;
    import udp_echo_app_stats_pkg::*;
    import beehive_udp_app_logger_msg::*;

`endif
