`ifndef NOC_DATACTRL_CONVERT_SVH
`define NOC_DATACTRL_CONVERT_SVH
    `include "noc_defs.vh"
    import beehive_noc_msg::*;
    import beehive_ctrl_noc_msg::*;

`endif
