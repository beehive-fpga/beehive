`ifndef ECHO_APP_STATS_DEFS_SVH
`define ECHO_APP_STATS_DEFS_SVH
    import echo_app_stats_pkg::*;

    import beehive_echo_app_logger_msg::*;

`endif
