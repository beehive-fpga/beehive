`ifndef MASKED_MEM_DEFS_SVH
`define MASKED_MEM_DEFS_SVH
    `include "noc_defs.vh"

    import beehive_noc_msg::*;

`endif
