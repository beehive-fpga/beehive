`ifndef ETH_TX_TILE_DEFS
`define ETH_TX_TILE_DEFS
    
    import beehive_eth_msg::*;
    import beehive_noc_msg::*;

    import packet_struct_pkg::*;
    
    `include "packet_defs.vh"    
    `include "noc_defs.vh"
    `include "soc_defs.vh"
`endif
