`ifndef MRP_TX_DEFS_SVH
`define MRP_TX_DEFS_SVH
    `include "noc_defs.vh"
    `include "noc_struct_defs.vh"
    `include "soc_defs.vh"
    `include "packet_defs.vh"
    
    import beehive_udp_msg::*;
    import beehive_noc_msg::*;
    import mrp_tx_pkg::*;
    import beehive_topology::*;

`endif
