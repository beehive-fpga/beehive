`ifndef SIMPLE_LOG_UDP_NOC_READ_DEFS
`define SIMPLE_LOG_UDP_NOC_READ_DEFS

    import beehive_topology::*;
    import beehive_noc_msg::*;
    import beehive_udp_msg::*;
    import simple_log_udp_noc_read_pkg::*;
    `include "noc_defs.vh"
`endif
