`ifndef TCP_LOGGER_READ_DEFS_SVH
`define TCP_LOGGER_READ_DEFS_SVH
    `include "noc_defs.vh"

    import beehive_noc_msg::*;
    import beehive_udp_msg::*;
    import beehive_topology::*;

    import tcp_logger_pkg::*;
`endif
