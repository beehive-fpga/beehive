`ifndef UDP_ECHO_APP_DEFS_SVH
`define UDP_ECHO_APP_DEFS_SVH
    import udp_echo_app_pkg::*;
    import beehive_topology::*;
    import beehive_noc_msg::*;
    import beehive_udp_msg::*;

    `include "noc_defs.vh"
    `include "packet_defs.vh"

`endif
