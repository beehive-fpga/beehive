`ifndef BEEHIVE_TCP_ENGINE_DEFS
`define BEEHIVE_TCP_ENGINE_DEFS
    `include "packet_defs.vh"
    `include "soc_defs.vh"

    import packet_struct_pkg::*;
    import tcp_pkg::*;
    import tcp_misc_pkg::*;
`endif
