`ifndef MRP_DEFS_SVH
`define MRP_DEFS_SVH

`include "packet_defs.vh"
`include "soc_defs.vh"

import mrp_pkg::*;

`endif
