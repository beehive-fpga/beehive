`ifndef NOC_ROUTER_BLOCK_DEFS_SVH
`define NOC_ROUTER_BLOCK_DEFS_SVH
    `include "noc_defs.vh"

`endif
