package beehive_topology;
    localparam UDP_TX_TILE_X = 1;
    localparam UDP_TX_TILE_Y = 1;
    localparam PKT_IF_FBITS = 9;

    localparam APP_SETUP_PORT = 52001;
    localparam APP_PORT = 52000;
endpackage
