`ifndef TCP_MSG_POLLER_DEFS_SVH
`define TCP_MSG_POLLER_DEFS_SVH
    `include "noc_defs.vh"

    import tcp_msg_poller_pkg::*;
    import tcp_pkg::*;
`endif
