`ifndef IP_REWRITE_NOC_PIPE_DEFS_SVH
`define IP_REWRITE_NOC_PIPE_DEFS_SVH
    import ip_rewrite_noc_pipe_pkg::*;
    import beehive_ip_msg::*;
    import beehive_noc_msg::*;
    
    `include "packet_defs.vh"
    `include "noc_defs.vh"

`endif
