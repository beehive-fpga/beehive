`ifndef IP_ENCAP_TX_DEFS
`define IP_ENCAP_TX_DEFS
    `include "packet_defs.vh"
    `include "noc_defs.vh"
    `include "noc_struct_defs.vh" 
    `include "bsg_defines.v"

    import ip_encap_tx_pkg::*;
    import beehive_ip_msg::*;
    import beehive_topology::*;
`endif

