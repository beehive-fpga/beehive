`ifndef LOGGER_TILE_DEFS
`define LOGGER_TILE_DEFS
    `include "noc_defs.vh"

    import beehive_noc_msg::*;
    import beehive_tcp_logger_msg::*;
    import tcp_logger_pkg::*;
`endif
