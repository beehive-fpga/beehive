package eth_tx_tile_pkg;
    
endpackage 
