`ifndef TO_IP_DEFS_SVH
`define TO_IP_DEFS_SVH
    `include "noc_defs.vh"
    `include "soc_defs.vh"
    `include "packet_defs.vh"

    import beehive_noc_msg::*;
    import beehive_ip_msg::*;
    import beehive_topology::*;
    import to_ip_tx_pkg::*;
`endif
