`ifndef RS_ENCODE_STATS_DEFS_SVH
`define RS_ENCODE_STATS_DEFS_SVH

    import rs_encode_stats_pkg::*; 

    `include "noc_defs.vh"

`endif
