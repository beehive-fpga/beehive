package ip_encap_tx_pkg;

    localparam IP_CAM_ELS = 8;
    localparam IP_CAM_INIT_ELS = 2;
endpackage
