`ifndef ECHO_APP_DEFS_SVH
`define ECHO_APP_DEFS_SVH

    `include "noc_defs.vh"

    import echo_app_pkg::*;
    import beehive_noc_msg::*;
    import beehive_tcp_msg::*;
    import beehive_topology::*;

    import tcp_pkg::*;
`endif
