`ifndef INGRESS_LOAD_BALANCE_DEFS_SVH
`define INGRESS_LOAD_BALANCE_DEFS_SVH

    `include "noc_defs.vh"
    `include "soc_defs.vh"

`endif
