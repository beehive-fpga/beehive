module demux_one_hot #(
     parameter NUM_OUTPUTS = -1
    ,parameter INPUT_WIDTH = -1
)(
     input  logic   [NUM_OUTPUTS-1:0]                    input_sel
    ,input  logic                    [INPUT_WIDTH-1:0]   data_input
    ,output logic   [NUM_OUTPUTS-1:0][INPUT_WIDTH-1:0]   data_outputs
);

    genvar i;
    generate
        for (i = 0; i < NUM_OUTPUTS; i = i + 1) begin
            always_comb begin
                data_outputs[i] = {(INPUT_WIDTH){input_sel[i]}} & data_input;
            end
        end
    endgenerate
endmodule
