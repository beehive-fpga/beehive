`ifndef ETH_LATENCY_STATS_DEFS
`define ETH_LATENCY_STATS_DEFS

    import beehive_noc_msg::*;
    import beehive_udp_msg::*;
    import beehive_eth_latency_logger_msg::*;
    import eth_latency_stats_pkg::*;

    `include "noc_defs.vh"

`endif
