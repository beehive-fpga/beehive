`ifndef RR_SCHEDULER_DEFS
`define RR_SCHEDULER_DEFS

    `include "noc_defs.vh"
    import scheduler_pkg::*;
    import beehive_noc_msg::*;

`endif
