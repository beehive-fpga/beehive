`ifndef TCP_LOGGER_RECORD_DEFS_SVH
`define TCP_LOGGER_RECORD_DEFS_SVH
    `include "noc_defs.vh"
    import packet_struct_pkg::*;

    import tcp_logger_pkg::*;
    import beehive_noc_msg::*;
    import beehive_ip_msg::*;
    import beehive_topology::*;

`endif
