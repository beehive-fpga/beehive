package rr_scheduler_pkg;
endpackage
