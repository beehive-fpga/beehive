`ifndef IP_REWRITE_MANAGER_DEFS_SVH
`define IP_REWRITE_MANAGER_DEFS_SVH
    `include "noc_defs.vh"
   
    import ip_rewrite_manager_pkg::*;

    import beehive_ip_rewrite_msg::*;
    import beehive_noc_msg::*;
    import beehive_tcp_msg::*;

`endif
