`ifndef UDP_TX_TILE_DEFS
`define UDP_TX_TILE_DEFS

    `include "noc_defs.vh"
    `include "packet_defs.vh"

    import packet_struct_pkg::*;

    import beehive_udp_msg::*;
    import beehive_ip_msg::*;
    import beehive_noc_msg::*;
    import udp_tx_tile_pkg::*;
    import beehive_topology::*;

`endif
